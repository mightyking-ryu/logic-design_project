`timescale 1ns/1ps

module pseudo_random(input  clk, rstn, gen, input [31:0] N, output [31:0] q, output gen_end);
    //Implement pseudo random number generator
    
    
     
endmodule
