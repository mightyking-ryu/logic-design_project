module unpack_mod(
    input clk,rstn,sel_bit,gen,
    input [31:0] message0,message1,N,
    input [31:0] rand_val,
    output [31:0] unpack_res,
    output gen_end
    );

    //Implement unpack_mod module
    //This module calculates 
    //m_b = (m_b' -k) mod N
    //on receiver side

    
       
endmodule
